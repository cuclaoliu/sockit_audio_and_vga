// nios_core.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module nios_core (
		output wire        audio_xck,                                  //            audio.xck
		input  wire        audio_daclrc,                               //                 .daclrc
		output wire        audio_dacdat,                               //                 .dacdat
		input  wire        audio_bclk,                                 //                 .bclk
		input  wire        audio_adclrc,                               //                 .adclrc
		input  wire        audio_adcdat,                               //                 .adcdat
		input  wire        clk_clk,                                    //              clk.clk
		input  wire        ddr3_pll_ref_clk_clk,                       // ddr3_pll_ref_clk.clk
		output wire        ddr3_pll_sharing_pll_mem_clk,               // ddr3_pll_sharing.pll_mem_clk
		output wire        ddr3_pll_sharing_pll_write_clk,             //                 .pll_write_clk
		output wire        ddr3_pll_sharing_pll_locked,                //                 .pll_locked
		output wire        ddr3_pll_sharing_pll_write_clk_pre_phy_clk, //                 .pll_write_clk_pre_phy_clk
		output wire        ddr3_pll_sharing_pll_addr_cmd_clk,          //                 .pll_addr_cmd_clk
		output wire        ddr3_pll_sharing_pll_avl_clk,               //                 .pll_avl_clk
		output wire        ddr3_pll_sharing_pll_config_clk,            //                 .pll_config_clk
		output wire        ddr3_pll_sharing_pll_mem_phy_clk,           //                 .pll_mem_phy_clk
		output wire        ddr3_pll_sharing_afi_phy_clk,               //                 .afi_phy_clk
		output wire        ddr3_pll_sharing_pll_avl_phy_clk,           //                 .pll_avl_phy_clk
		output wire        ddr3_status_local_init_done,                //      ddr3_status.local_init_done
		output wire        ddr3_status_local_cal_success,              //                 .local_cal_success
		output wire        ddr3_status_local_cal_fail,                 //                 .local_cal_fail
		output wire        i2c_scl_export,                             //          i2c_scl.export
		inout  wire        i2c_sda_export,                             //          i2c_sda.export
		output wire [14:0] memory_mem_a,                               //           memory.mem_a
		output wire [2:0]  memory_mem_ba,                              //                 .mem_ba
		output wire [0:0]  memory_mem_ck,                              //                 .mem_ck
		output wire [0:0]  memory_mem_ck_n,                            //                 .mem_ck_n
		output wire [0:0]  memory_mem_cke,                             //                 .mem_cke
		output wire [0:0]  memory_mem_cs_n,                            //                 .mem_cs_n
		output wire [3:0]  memory_mem_dm,                              //                 .mem_dm
		output wire [0:0]  memory_mem_ras_n,                           //                 .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                           //                 .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                            //                 .mem_we_n
		output wire        memory_mem_reset_n,                         //                 .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                              //                 .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                             //                 .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                           //                 .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                             //                 .mem_odt
		input  wire        oct_rzqin,                                  //              oct.rzqin
		input  wire [3:0]  pio_key_export,                             //          pio_key.export
		output wire [3:0]  pio_led_export,                             //          pio_led.export
		input  wire [3:0]  pio_sw_export,                              //           pio_sw.export
		input  wire        reset_reset_n,                              //            reset.reset_n
		output wire        vga_vga_hs,                                 //              vga.vga_hs
		output wire        vga_vga_vs,                                 //                 .vga_vs
		output wire        vga_vga_de,                                 //                 .vga_de
		output wire [7:0]  vga_vga_r,                                  //                 .vga_r
		output wire [7:0]  vga_vga_g,                                  //                 .vga_g
		output wire [7:0]  vga_vga_b,                                  //                 .vga_b
		output wire        vga_clk_clk                                 //          vga_clk.clk
	);

	wire          pll_sys_outclk0_clk;                                       // pll_sys:outclk_0 -> [cpu:clk, cpu_peripheral_bridge:s0_clk, data_buffer:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_sys_outclk0_clk, onchip_memory:clk, rst_controller_001:clk, sysid_qsys:clock, timer:clk]
	wire          pll_audio_outclk0_clk;                                     // pll_audio:outclk_0 -> [audio:avs_s1_clk, mm_interconnect_0:pll_audio_outclk0_clk, rst_controller:clk]
	wire          pll_sys_outclk1_clk;                                       // pll_sys:outclk_1 -> [cpu_peripheral_bridge:m0_clk, i2c_scl:clk, i2c_sda:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mm_interconnect_1:pll_sys_outclk1_clk, pio_key:clk, pio_led:clk, pio_sw:clk, rst_controller_002:clk]
	wire   [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire          cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire          cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [28:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire    [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire          cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire          cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire          cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire   [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire   [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire   [28:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire          cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire          cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [15:0] mm_interconnect_0_audio_avalon_slave_readdata;             // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire    [2:0] mm_interconnect_0_audio_avalon_slave_address;              // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire          mm_interconnect_0_audio_avalon_slave_read;                 // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire          mm_interconnect_0_audio_avalon_slave_write;                // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire   [15:0] mm_interconnect_0_audio_avalon_slave_writedata;            // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire          mm_interconnect_0_vpg_avalon_slave_chipselect;             // mm_interconnect_0:vpg_avalon_slave_chipselect -> vpg:avalon_slave_cs_n
	wire    [7:0] mm_interconnect_0_vpg_avalon_slave_readdata;               // vpg:avalon_slave_readdata -> mm_interconnect_0:vpg_avalon_slave_readdata
	wire          mm_interconnect_0_vpg_avalon_slave_read;                   // mm_interconnect_0:vpg_avalon_slave_read -> vpg:avalon_slave_read
	wire          mm_interconnect_0_vpg_avalon_slave_write;                  // mm_interconnect_0:vpg_avalon_slave_write -> vpg:avalon_slave_write
	wire    [7:0] mm_interconnect_0_vpg_avalon_slave_writedata;              // mm_interconnect_0:vpg_avalon_slave_writedata -> vpg:avalon_slave_writedata
	wire          mm_interconnect_0_ddr3_avl_beginbursttransfer;             // mm_interconnect_0:ddr3_avl_beginbursttransfer -> ddr3:avl_burstbegin
	wire  [127:0] mm_interconnect_0_ddr3_avl_readdata;                       // ddr3:avl_rdata -> mm_interconnect_0:ddr3_avl_readdata
	wire          mm_interconnect_0_ddr3_avl_waitrequest;                    // ddr3:avl_ready -> mm_interconnect_0:ddr3_avl_waitrequest
	wire   [23:0] mm_interconnect_0_ddr3_avl_address;                        // mm_interconnect_0:ddr3_avl_address -> ddr3:avl_addr
	wire          mm_interconnect_0_ddr3_avl_read;                           // mm_interconnect_0:ddr3_avl_read -> ddr3:avl_read_req
	wire   [15:0] mm_interconnect_0_ddr3_avl_byteenable;                     // mm_interconnect_0:ddr3_avl_byteenable -> ddr3:avl_be
	wire          mm_interconnect_0_ddr3_avl_readdatavalid;                  // ddr3:avl_rdata_valid -> mm_interconnect_0:ddr3_avl_readdatavalid
	wire          mm_interconnect_0_ddr3_avl_write;                          // mm_interconnect_0:ddr3_avl_write -> ddr3:avl_write_req
	wire  [127:0] mm_interconnect_0_ddr3_avl_writedata;                      // mm_interconnect_0:ddr3_avl_writedata -> ddr3:avl_wdata
	wire    [5:0] mm_interconnect_0_ddr3_avl_burstcount;                     // mm_interconnect_0:ddr3_avl_burstcount -> ddr3:avl_size
	wire          ddr3_afi_clk_clk;                                          // ddr3:afi_clk -> [mm_interconnect_0:ddr3_afi_clk_clk, rst_controller_009:clk]
	wire   [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire          mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire          mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire          mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_0_cpu_peripheral_bridge_s0_readdata;       // cpu_peripheral_bridge:s0_readdata -> mm_interconnect_0:cpu_peripheral_bridge_s0_readdata
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest;    // cpu_peripheral_bridge:s0_waitrequest -> mm_interconnect_0:cpu_peripheral_bridge_s0_waitrequest
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess;    // mm_interconnect_0:cpu_peripheral_bridge_s0_debugaccess -> cpu_peripheral_bridge:s0_debugaccess
	wire    [8:0] mm_interconnect_0_cpu_peripheral_bridge_s0_address;        // mm_interconnect_0:cpu_peripheral_bridge_s0_address -> cpu_peripheral_bridge:s0_address
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_read;           // mm_interconnect_0:cpu_peripheral_bridge_s0_read -> cpu_peripheral_bridge:s0_read
	wire    [3:0] mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable;     // mm_interconnect_0:cpu_peripheral_bridge_s0_byteenable -> cpu_peripheral_bridge:s0_byteenable
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid;  // cpu_peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:cpu_peripheral_bridge_s0_readdatavalid
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_write;          // mm_interconnect_0:cpu_peripheral_bridge_s0_write -> cpu_peripheral_bridge:s0_write
	wire   [31:0] mm_interconnect_0_cpu_peripheral_bridge_s0_writedata;      // mm_interconnect_0:cpu_peripheral_bridge_s0_writedata -> cpu_peripheral_bridge:s0_writedata
	wire    [0:0] mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount;     // mm_interconnect_0:cpu_peripheral_bridge_s0_burstcount -> cpu_peripheral_bridge:s0_burstcount
	wire          mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire   [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [15:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire    [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire          mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire   [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire          mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire          mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire   [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire    [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire          mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire   [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire          mm_interconnect_0_data_buffer_s1_chipselect;               // mm_interconnect_0:data_buffer_s1_chipselect -> data_buffer:chipselect
	wire   [31:0] mm_interconnect_0_data_buffer_s1_readdata;                 // data_buffer:readdata -> mm_interconnect_0:data_buffer_s1_readdata
	wire    [9:0] mm_interconnect_0_data_buffer_s1_address;                  // mm_interconnect_0:data_buffer_s1_address -> data_buffer:address
	wire    [3:0] mm_interconnect_0_data_buffer_s1_byteenable;               // mm_interconnect_0:data_buffer_s1_byteenable -> data_buffer:byteenable
	wire          mm_interconnect_0_data_buffer_s1_write;                    // mm_interconnect_0:data_buffer_s1_write -> data_buffer:write
	wire   [31:0] mm_interconnect_0_data_buffer_s1_writedata;                // mm_interconnect_0:data_buffer_s1_writedata -> data_buffer:writedata
	wire          mm_interconnect_0_data_buffer_s1_clken;                    // mm_interconnect_0:data_buffer_s1_clken -> data_buffer:clken
	wire          cpu_peripheral_bridge_m0_waitrequest;                      // mm_interconnect_1:cpu_peripheral_bridge_m0_waitrequest -> cpu_peripheral_bridge:m0_waitrequest
	wire   [31:0] cpu_peripheral_bridge_m0_readdata;                         // mm_interconnect_1:cpu_peripheral_bridge_m0_readdata -> cpu_peripheral_bridge:m0_readdata
	wire          cpu_peripheral_bridge_m0_debugaccess;                      // cpu_peripheral_bridge:m0_debugaccess -> mm_interconnect_1:cpu_peripheral_bridge_m0_debugaccess
	wire    [8:0] cpu_peripheral_bridge_m0_address;                          // cpu_peripheral_bridge:m0_address -> mm_interconnect_1:cpu_peripheral_bridge_m0_address
	wire          cpu_peripheral_bridge_m0_read;                             // cpu_peripheral_bridge:m0_read -> mm_interconnect_1:cpu_peripheral_bridge_m0_read
	wire    [3:0] cpu_peripheral_bridge_m0_byteenable;                       // cpu_peripheral_bridge:m0_byteenable -> mm_interconnect_1:cpu_peripheral_bridge_m0_byteenable
	wire          cpu_peripheral_bridge_m0_readdatavalid;                    // mm_interconnect_1:cpu_peripheral_bridge_m0_readdatavalid -> cpu_peripheral_bridge:m0_readdatavalid
	wire   [31:0] cpu_peripheral_bridge_m0_writedata;                        // cpu_peripheral_bridge:m0_writedata -> mm_interconnect_1:cpu_peripheral_bridge_m0_writedata
	wire          cpu_peripheral_bridge_m0_write;                            // cpu_peripheral_bridge:m0_write -> mm_interconnect_1:cpu_peripheral_bridge_m0_write
	wire    [0:0] cpu_peripheral_bridge_m0_burstcount;                       // cpu_peripheral_bridge:m0_burstcount -> mm_interconnect_1:cpu_peripheral_bridge_m0_burstcount
	wire          mm_interconnect_1_pio_key_s1_chipselect;                   // mm_interconnect_1:pio_key_s1_chipselect -> pio_key:chipselect
	wire   [31:0] mm_interconnect_1_pio_key_s1_readdata;                     // pio_key:readdata -> mm_interconnect_1:pio_key_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_key_s1_address;                      // mm_interconnect_1:pio_key_s1_address -> pio_key:address
	wire          mm_interconnect_1_pio_key_s1_write;                        // mm_interconnect_1:pio_key_s1_write -> pio_key:write_n
	wire   [31:0] mm_interconnect_1_pio_key_s1_writedata;                    // mm_interconnect_1:pio_key_s1_writedata -> pio_key:writedata
	wire          mm_interconnect_1_pio_led_s1_chipselect;                   // mm_interconnect_1:pio_led_s1_chipselect -> pio_led:chipselect
	wire   [31:0] mm_interconnect_1_pio_led_s1_readdata;                     // pio_led:readdata -> mm_interconnect_1:pio_led_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_led_s1_address;                      // mm_interconnect_1:pio_led_s1_address -> pio_led:address
	wire          mm_interconnect_1_pio_led_s1_write;                        // mm_interconnect_1:pio_led_s1_write -> pio_led:write_n
	wire   [31:0] mm_interconnect_1_pio_led_s1_writedata;                    // mm_interconnect_1:pio_led_s1_writedata -> pio_led:writedata
	wire          mm_interconnect_1_pio_sw_s1_chipselect;                    // mm_interconnect_1:pio_sw_s1_chipselect -> pio_sw:chipselect
	wire   [31:0] mm_interconnect_1_pio_sw_s1_readdata;                      // pio_sw:readdata -> mm_interconnect_1:pio_sw_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_sw_s1_address;                       // mm_interconnect_1:pio_sw_s1_address -> pio_sw:address
	wire          mm_interconnect_1_pio_sw_s1_write;                         // mm_interconnect_1:pio_sw_s1_write -> pio_sw:write_n
	wire   [31:0] mm_interconnect_1_pio_sw_s1_writedata;                     // mm_interconnect_1:pio_sw_s1_writedata -> pio_sw:writedata
	wire          mm_interconnect_1_i2c_scl_s1_chipselect;                   // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire   [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                     // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire    [1:0] mm_interconnect_1_i2c_scl_s1_address;                      // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire          mm_interconnect_1_i2c_scl_s1_write;                        // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire   [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                    // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire          mm_interconnect_1_i2c_sda_s1_chipselect;                   // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire   [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                     // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire    [1:0] mm_interconnect_1_i2c_sda_s1_address;                      // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire          mm_interconnect_1_i2c_sda_s1_write;                        // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire   [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                    // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire          irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver3_irq;                                  // timer:irq -> irq_mapper:receiver3_irq
	wire   [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire          irq_mapper_receiver1_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                             // pio_key:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver2_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                         // pio_sw:irq -> irq_synchronizer_001:receiver_irq
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [audio:avs_s1_reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset]
	wire          ddr3_afi_reset_reset;                                      // ddr3:afi_reset_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0, rst_controller_007:reset_in0, rst_controller_008:reset_in0]
	wire          ddr3_afi_reset_export_reset;                               // ddr3:afi_reset_export_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_005:reset_in1, rst_controller_006:reset_in1, rst_controller_007:reset_in1, rst_controller_008:reset_in1]
	wire          cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller:reset_in3, rst_controller_001:reset_in3, rst_controller_002:reset_in3, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in3, rst_controller_006:reset_in3, rst_controller_007:reset_in3, rst_controller_008:reset_in3, rst_controller_009:reset_in1]
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [cpu:reset_n, cpu_peripheral_bridge:s0_reset, data_buffer:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset, sysid_qsys:reset_n, timer:reset_n]
	wire          rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [cpu:reset_req, data_buffer:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [cpu_peripheral_bridge:m0_reset, i2c_scl:reset_n, i2c_sda:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_1:cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset_reset, pio_key:reset_n, pio_led:reset_n, pio_sw:reset_n]
	wire          rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> ddr3:global_reset_n
	wire          rst_controller_004_reset_out_reset;                        // rst_controller_004:reset_out -> ddr3:soft_reset_n
	wire          rst_controller_005_reset_out_reset;                        // rst_controller_005:reset_out -> pll_audio:rst
	wire          rst_controller_006_reset_out_reset;                        // rst_controller_006:reset_out -> pll_sys:rst
	wire          rst_controller_007_reset_out_reset;                        // rst_controller_007:reset_out -> vga_pll:rst
	wire          rst_controller_008_reset_out_reset;                        // rst_controller_008:reset_out -> [mm_interconnect_0:vpg_reset_reset_bridge_in_reset_reset, vpg:reset_n]
	wire          rst_controller_009_reset_out_reset;                        // rst_controller_009:reset_out -> [mm_interconnect_0:ddr3_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ddr3_soft_reset_reset_bridge_in_reset_reset]

	AUDIO_IF audio (
		.avs_s1_address   (mm_interconnect_0_audio_avalon_slave_address),   // avalon_slave.address
		.avs_s1_read      (mm_interconnect_0_audio_avalon_slave_read),      //             .read
		.avs_s1_readdata  (mm_interconnect_0_audio_avalon_slave_readdata),  //             .readdata
		.avs_s1_write     (mm_interconnect_0_audio_avalon_slave_write),     //             .write
		.avs_s1_writedata (mm_interconnect_0_audio_avalon_slave_writedata), //             .writedata
		.avs_s1_clk       (pll_audio_outclk0_clk),                          //        clock.clk
		.avs_s1_reset     (rst_controller_reset_out_reset),                 //        reset.reset
		.audio_XCK        (audio_xck),                                      //      conduit.xck
		.audio_DACLRC     (audio_daclrc),                                   //             .daclrc
		.audio_DACDAT     (audio_dacdat),                                   //             .dacdat
		.audio_BCLK       (audio_bclk),                                     //             .bclk
		.audio_ADCLRC     (audio_adclrc),                                   //             .adclrc
		.audio_ADCDAT     (audio_adcdat)                                    //             .adcdat
	);

	nios_core_cpu cpu (
		.clk                                 (pll_sys_outclk0_clk),                               //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_peripheral_bridge (
		.m0_clk           (pll_sys_outclk1_clk),                                      //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (pll_sys_outclk0_clk),                                      //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cpu_peripheral_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_cpu_peripheral_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_cpu_peripheral_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_cpu_peripheral_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_cpu_peripheral_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_peripheral_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (cpu_peripheral_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (cpu_peripheral_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (cpu_peripheral_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (cpu_peripheral_bridge_m0_writedata),                       //         .writedata
		.m0_address       (cpu_peripheral_bridge_m0_address),                         //         .address
		.m0_write         (cpu_peripheral_bridge_m0_write),                           //         .write
		.m0_read          (cpu_peripheral_bridge_m0_read),                            //         .read
		.m0_byteenable    (cpu_peripheral_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (cpu_peripheral_bridge_m0_debugaccess)                      //         .debugaccess
	);

	nios_core_data_buffer data_buffer (
		.clk        (pll_sys_outclk0_clk),                         //   clk1.clk
		.address    (mm_interconnect_0_data_buffer_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_buffer_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_buffer_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_buffer_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_buffer_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_buffer_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_buffer_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	nios_core_ddr3 ddr3 (
		.pll_ref_clk               (ddr3_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n            (~rst_controller_003_reset_out_reset),           //     global_reset.reset_n
		.soft_reset_n              (~rst_controller_004_reset_out_reset),           //       soft_reset.reset_n
		.afi_clk                   (ddr3_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                              //     afi_half_clk.clk
		.afi_reset_n               (ddr3_afi_reset_reset),                          //        afi_reset.reset_n
		.afi_reset_export_n        (ddr3_afi_reset_export_reset),                   // afi_reset_export.reset_n
		.mem_a                     (memory_mem_a),                                  //           memory.mem_a
		.mem_ba                    (memory_mem_ba),                                 //                 .mem_ba
		.mem_ck                    (memory_mem_ck),                                 //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                               //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                               //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                                 //                 .mem_dm
		.mem_ras_n                 (memory_mem_ras_n),                              //                 .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                              //                 .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                               //                 .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                            //                 .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                 //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                              //                 .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                //                 .mem_odt
		.avl_ready                 (mm_interconnect_0_ddr3_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_0_ddr3_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_0_ddr3_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_0_ddr3_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_0_ddr3_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_0_ddr3_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_0_ddr3_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_0_ddr3_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_0_ddr3_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_0_ddr3_avl_burstcount),         //                 .burstcount
		.local_init_done           (ddr3_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (ddr3_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (ddr3_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                                     //              oct.rzqin
		.pll_mem_clk               (ddr3_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk             (ddr3_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked                (ddr3_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_write_clk_pre_phy_clk (ddr3_pll_sharing_pll_write_clk_pre_phy_clk),    //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (ddr3_pll_sharing_pll_addr_cmd_clk),             //                 .pll_addr_cmd_clk
		.pll_avl_clk               (ddr3_pll_sharing_pll_avl_clk),                  //                 .pll_avl_clk
		.pll_config_clk            (ddr3_pll_sharing_pll_config_clk),               //                 .pll_config_clk
		.pll_mem_phy_clk           (ddr3_pll_sharing_pll_mem_phy_clk),              //                 .pll_mem_phy_clk
		.afi_phy_clk               (ddr3_pll_sharing_afi_phy_clk),                  //                 .afi_phy_clk
		.pll_avl_phy_clk           (ddr3_pll_sharing_pll_avl_phy_clk)               //                 .pll_avl_phy_clk
	);

	nios_core_i2c_scl i2c_scl (
		.clk        (pll_sys_outclk1_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_export)                           // external_connection.export
	);

	nios_core_i2c_sda i2c_sda (
		.clk        (pll_sys_outclk1_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_export)                           // external_connection.export
	);

	nios_core_jtag_uart jtag_uart (
		.clk            (pll_sys_outclk0_clk),                                       //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios_core_onchip_memory onchip_memory (
		.clk        (pll_sys_outclk0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	nios_core_pio_key pio_key (
		.clk        (pll_sys_outclk1_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_pio_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_key_s1_readdata),   //                    .readdata
		.in_port    (pio_key_export),                          // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)            //                 irq.irq
	);

	nios_core_pio_led pio_led (
		.clk        (pll_sys_outclk1_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	nios_core_pio_key pio_sw (
		.clk        (pll_sys_outclk1_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_pio_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_sw_s1_readdata),   //                    .readdata
		.in_port    (pio_sw_export),                          // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)       //                 irq.irq
	);

	nios_core_pll_audio pll_audio (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_005_reset_out_reset), //   reset.reset
		.outclk_0 (pll_audio_outclk0_clk),              // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	nios_core_pll_sys pll_sys (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_006_reset_out_reset), //   reset.reset
		.outclk_0 (pll_sys_outclk0_clk),                // outclk0.clk
		.outclk_1 (pll_sys_outclk1_clk),                // outclk1.clk
		.locked   ()                                    // (terminated)
	);

	nios_core_sysid_qsys sysid_qsys (
		.clock    (pll_sys_outclk0_clk),                                 //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	nios_core_timer timer (
		.clk        (pll_sys_outclk0_clk),                   //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
	);

	nios_core_vga_pll vga_pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_007_reset_out_reset), //   reset.reset
		.outclk_0 (vga_clk_clk),                        // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	vpg #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (24),
		.READY_LATENCY    (0),
		.MAX_CHANNEL      (0),
		.H_DISP           (640),
		.H_FPORCH         (16),
		.H_SYNC           (96),
		.H_BPORCH         (48),
		.V_DISP           (480),
		.V_FPORCH         (10),
		.V_SYNC           (2),
		.V_BPORCH         (33)
	) vpg (
		.clk                    (vga_clk_clk),                                    //        clock.clk
		.reset_n                (~rst_controller_008_reset_out_reset),            //        reset.reset_n
		.vga_hs                 (vga_vga_hs),                                     //  conduit_end.vga_hs
		.vga_vs                 (vga_vga_vs),                                     //             .vga_vs
		.vga_de                 (vga_vga_de),                                     //             .vga_de
		.vga_r                  (vga_vga_r),                                      //             .vga_r
		.vga_g                  (vga_vga_g),                                      //             .vga_g
		.vga_b                  (vga_vga_b),                                      //             .vga_b
		.avalon_slave_write     (mm_interconnect_0_vpg_avalon_slave_write),       // avalon_slave.write
		.avalon_slave_writedata (mm_interconnect_0_vpg_avalon_slave_writedata),   //             .writedata
		.avalon_slave_read      (mm_interconnect_0_vpg_avalon_slave_read),        //             .read
		.avalon_slave_readdata  (mm_interconnect_0_vpg_avalon_slave_readdata),    //             .readdata
		.avalon_slave_cs_n      (~mm_interconnect_0_vpg_avalon_slave_chipselect)  //             .chipselect_n
	);

	nios_core_mm_interconnect_0 mm_interconnect_0 (
		.ddr3_afi_clk_clk                                      (ddr3_afi_clk_clk),                                          //                                    ddr3_afi_clk.clk
		.pll_audio_outclk0_clk                                 (pll_audio_outclk0_clk),                                     //                               pll_audio_outclk0.clk
		.pll_sys_outclk0_clk                                   (pll_sys_outclk0_clk),                                       //                                 pll_sys_outclk0.clk
		.vga_pll_outclk0_clk                                   (vga_clk_clk),                                               //                                 vga_pll_outclk0.clk
		.audio_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                            //               audio_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                 (rst_controller_001_reset_out_reset),                        //                 cpu_reset_reset_bridge_in_reset.reset
		.ddr3_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_009_reset_out_reset),                        // ddr3_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr3_soft_reset_reset_bridge_in_reset_reset           (rst_controller_009_reset_out_reset),                        //           ddr3_soft_reset_reset_bridge_in_reset.reset
		.vpg_reset_reset_bridge_in_reset_reset                 (rst_controller_008_reset_out_reset),                        //                 vpg_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                   //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                      //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                  //                                                .readdata
		.cpu_data_master_readdatavalid                         (cpu_data_master_readdatavalid),                             //                                                .readdatavalid
		.cpu_data_master_write                                 (cpu_data_master_write),                                     //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                 //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                            //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                               //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                           //                                                .readdata
		.cpu_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                      //                                                .readdatavalid
		.audio_avalon_slave_address                            (mm_interconnect_0_audio_avalon_slave_address),              //                              audio_avalon_slave.address
		.audio_avalon_slave_write                              (mm_interconnect_0_audio_avalon_slave_write),                //                                                .write
		.audio_avalon_slave_read                               (mm_interconnect_0_audio_avalon_slave_read),                 //                                                .read
		.audio_avalon_slave_readdata                           (mm_interconnect_0_audio_avalon_slave_readdata),             //                                                .readdata
		.audio_avalon_slave_writedata                          (mm_interconnect_0_audio_avalon_slave_writedata),            //                                                .writedata
		.cpu_debug_mem_slave_address                           (mm_interconnect_0_cpu_debug_mem_slave_address),             //                             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                             (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                                .write
		.cpu_debug_mem_slave_read                              (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                                .read
		.cpu_debug_mem_slave_readdata                          (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                                .readdata
		.cpu_debug_mem_slave_writedata                         (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                                .writedata
		.cpu_debug_mem_slave_byteenable                        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                                .byteenable
		.cpu_debug_mem_slave_waitrequest                       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                                .waitrequest
		.cpu_debug_mem_slave_debugaccess                       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                                .debugaccess
		.cpu_peripheral_bridge_s0_address                      (mm_interconnect_0_cpu_peripheral_bridge_s0_address),        //                        cpu_peripheral_bridge_s0.address
		.cpu_peripheral_bridge_s0_write                        (mm_interconnect_0_cpu_peripheral_bridge_s0_write),          //                                                .write
		.cpu_peripheral_bridge_s0_read                         (mm_interconnect_0_cpu_peripheral_bridge_s0_read),           //                                                .read
		.cpu_peripheral_bridge_s0_readdata                     (mm_interconnect_0_cpu_peripheral_bridge_s0_readdata),       //                                                .readdata
		.cpu_peripheral_bridge_s0_writedata                    (mm_interconnect_0_cpu_peripheral_bridge_s0_writedata),      //                                                .writedata
		.cpu_peripheral_bridge_s0_burstcount                   (mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount),     //                                                .burstcount
		.cpu_peripheral_bridge_s0_byteenable                   (mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable),     //                                                .byteenable
		.cpu_peripheral_bridge_s0_readdatavalid                (mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid),  //                                                .readdatavalid
		.cpu_peripheral_bridge_s0_waitrequest                  (mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest),    //                                                .waitrequest
		.cpu_peripheral_bridge_s0_debugaccess                  (mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess),    //                                                .debugaccess
		.data_buffer_s1_address                                (mm_interconnect_0_data_buffer_s1_address),                  //                                  data_buffer_s1.address
		.data_buffer_s1_write                                  (mm_interconnect_0_data_buffer_s1_write),                    //                                                .write
		.data_buffer_s1_readdata                               (mm_interconnect_0_data_buffer_s1_readdata),                 //                                                .readdata
		.data_buffer_s1_writedata                              (mm_interconnect_0_data_buffer_s1_writedata),                //                                                .writedata
		.data_buffer_s1_byteenable                             (mm_interconnect_0_data_buffer_s1_byteenable),               //                                                .byteenable
		.data_buffer_s1_chipselect                             (mm_interconnect_0_data_buffer_s1_chipselect),               //                                                .chipselect
		.data_buffer_s1_clken                                  (mm_interconnect_0_data_buffer_s1_clken),                    //                                                .clken
		.ddr3_avl_address                                      (mm_interconnect_0_ddr3_avl_address),                        //                                        ddr3_avl.address
		.ddr3_avl_write                                        (mm_interconnect_0_ddr3_avl_write),                          //                                                .write
		.ddr3_avl_read                                         (mm_interconnect_0_ddr3_avl_read),                           //                                                .read
		.ddr3_avl_readdata                                     (mm_interconnect_0_ddr3_avl_readdata),                       //                                                .readdata
		.ddr3_avl_writedata                                    (mm_interconnect_0_ddr3_avl_writedata),                      //                                                .writedata
		.ddr3_avl_beginbursttransfer                           (mm_interconnect_0_ddr3_avl_beginbursttransfer),             //                                                .beginbursttransfer
		.ddr3_avl_burstcount                                   (mm_interconnect_0_ddr3_avl_burstcount),                     //                                                .burstcount
		.ddr3_avl_byteenable                                   (mm_interconnect_0_ddr3_avl_byteenable),                     //                                                .byteenable
		.ddr3_avl_readdatavalid                                (mm_interconnect_0_ddr3_avl_readdatavalid),                  //                                                .readdatavalid
		.ddr3_avl_waitrequest                                  (~mm_interconnect_0_ddr3_avl_waitrequest),                   //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.onchip_memory_s1_address                              (mm_interconnect_0_onchip_memory_s1_address),                //                                onchip_memory_s1.address
		.onchip_memory_s1_write                                (mm_interconnect_0_onchip_memory_s1_write),                  //                                                .write
		.onchip_memory_s1_readdata                             (mm_interconnect_0_onchip_memory_s1_readdata),               //                                                .readdata
		.onchip_memory_s1_writedata                            (mm_interconnect_0_onchip_memory_s1_writedata),              //                                                .writedata
		.onchip_memory_s1_byteenable                           (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                                .byteenable
		.onchip_memory_s1_chipselect                           (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                                .chipselect
		.onchip_memory_s1_clken                                (mm_interconnect_0_onchip_memory_s1_clken),                  //                                                .clken
		.sysid_qsys_control_slave_address                      (mm_interconnect_0_sysid_qsys_control_slave_address),        //                        sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                     (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                                .readdata
		.timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                        //                                        timer_s1.address
		.timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                          //                                                .write
		.timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                       //                                                .readdata
		.timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                      //                                                .writedata
		.timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                     //                                                .chipselect
		.vpg_avalon_slave_write                                (mm_interconnect_0_vpg_avalon_slave_write),                  //                                vpg_avalon_slave.write
		.vpg_avalon_slave_read                                 (mm_interconnect_0_vpg_avalon_slave_read),                   //                                                .read
		.vpg_avalon_slave_readdata                             (mm_interconnect_0_vpg_avalon_slave_readdata),               //                                                .readdata
		.vpg_avalon_slave_writedata                            (mm_interconnect_0_vpg_avalon_slave_writedata),              //                                                .writedata
		.vpg_avalon_slave_chipselect                           (mm_interconnect_0_vpg_avalon_slave_chipselect)              //                                                .chipselect
	);

	nios_core_mm_interconnect_1 mm_interconnect_1 (
		.pll_sys_outclk1_clk                                        (pll_sys_outclk1_clk),                     //                                      pll_sys_outclk1.clk
		.cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),      // cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset.reset
		.cpu_peripheral_bridge_m0_address                           (cpu_peripheral_bridge_m0_address),        //                             cpu_peripheral_bridge_m0.address
		.cpu_peripheral_bridge_m0_waitrequest                       (cpu_peripheral_bridge_m0_waitrequest),    //                                                     .waitrequest
		.cpu_peripheral_bridge_m0_burstcount                        (cpu_peripheral_bridge_m0_burstcount),     //                                                     .burstcount
		.cpu_peripheral_bridge_m0_byteenable                        (cpu_peripheral_bridge_m0_byteenable),     //                                                     .byteenable
		.cpu_peripheral_bridge_m0_read                              (cpu_peripheral_bridge_m0_read),           //                                                     .read
		.cpu_peripheral_bridge_m0_readdata                          (cpu_peripheral_bridge_m0_readdata),       //                                                     .readdata
		.cpu_peripheral_bridge_m0_readdatavalid                     (cpu_peripheral_bridge_m0_readdatavalid),  //                                                     .readdatavalid
		.cpu_peripheral_bridge_m0_write                             (cpu_peripheral_bridge_m0_write),          //                                                     .write
		.cpu_peripheral_bridge_m0_writedata                         (cpu_peripheral_bridge_m0_writedata),      //                                                     .writedata
		.cpu_peripheral_bridge_m0_debugaccess                       (cpu_peripheral_bridge_m0_debugaccess),    //                                                     .debugaccess
		.i2c_scl_s1_address                                         (mm_interconnect_1_i2c_scl_s1_address),    //                                           i2c_scl_s1.address
		.i2c_scl_s1_write                                           (mm_interconnect_1_i2c_scl_s1_write),      //                                                     .write
		.i2c_scl_s1_readdata                                        (mm_interconnect_1_i2c_scl_s1_readdata),   //                                                     .readdata
		.i2c_scl_s1_writedata                                       (mm_interconnect_1_i2c_scl_s1_writedata),  //                                                     .writedata
		.i2c_scl_s1_chipselect                                      (mm_interconnect_1_i2c_scl_s1_chipselect), //                                                     .chipselect
		.i2c_sda_s1_address                                         (mm_interconnect_1_i2c_sda_s1_address),    //                                           i2c_sda_s1.address
		.i2c_sda_s1_write                                           (mm_interconnect_1_i2c_sda_s1_write),      //                                                     .write
		.i2c_sda_s1_readdata                                        (mm_interconnect_1_i2c_sda_s1_readdata),   //                                                     .readdata
		.i2c_sda_s1_writedata                                       (mm_interconnect_1_i2c_sda_s1_writedata),  //                                                     .writedata
		.i2c_sda_s1_chipselect                                      (mm_interconnect_1_i2c_sda_s1_chipselect), //                                                     .chipselect
		.pio_key_s1_address                                         (mm_interconnect_1_pio_key_s1_address),    //                                           pio_key_s1.address
		.pio_key_s1_write                                           (mm_interconnect_1_pio_key_s1_write),      //                                                     .write
		.pio_key_s1_readdata                                        (mm_interconnect_1_pio_key_s1_readdata),   //                                                     .readdata
		.pio_key_s1_writedata                                       (mm_interconnect_1_pio_key_s1_writedata),  //                                                     .writedata
		.pio_key_s1_chipselect                                      (mm_interconnect_1_pio_key_s1_chipselect), //                                                     .chipselect
		.pio_led_s1_address                                         (mm_interconnect_1_pio_led_s1_address),    //                                           pio_led_s1.address
		.pio_led_s1_write                                           (mm_interconnect_1_pio_led_s1_write),      //                                                     .write
		.pio_led_s1_readdata                                        (mm_interconnect_1_pio_led_s1_readdata),   //                                                     .readdata
		.pio_led_s1_writedata                                       (mm_interconnect_1_pio_led_s1_writedata),  //                                                     .writedata
		.pio_led_s1_chipselect                                      (mm_interconnect_1_pio_led_s1_chipselect), //                                                     .chipselect
		.pio_sw_s1_address                                          (mm_interconnect_1_pio_sw_s1_address),     //                                            pio_sw_s1.address
		.pio_sw_s1_write                                            (mm_interconnect_1_pio_sw_s1_write),       //                                                     .write
		.pio_sw_s1_readdata                                         (mm_interconnect_1_pio_sw_s1_readdata),    //                                                     .readdata
		.pio_sw_s1_writedata                                        (mm_interconnect_1_pio_sw_s1_writedata),   //                                                     .writedata
		.pio_sw_s1_chipselect                                       (mm_interconnect_1_pio_sw_s1_chipselect)   //                                                     .chipselect
	);

	nios_core_irq_mapper irq_mapper (
		.clk           (pll_sys_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_sys_outclk1_clk),                //       receiver_clk.clk
		.sender_clk     (pll_sys_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_sys_outclk1_clk),                //       receiver_clk.clk
		.sender_clk     (pll_sys_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~ddr3_afi_reset_reset),          // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),   // reset_in1.reset
		.reset_in2      (~reset_reset_n),                 // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),  // reset_in3.reset
		.clk            (pll_audio_outclk0_clk),          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~ddr3_afi_reset_reset),                  // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),           // reset_in1.reset
		.reset_in2      (~reset_reset_n),                         // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),          // reset_in3.reset
		.clk            (pll_sys_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),       // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),      // reset_in3.reset
		.clk            (pll_sys_outclk1_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),       // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),      // reset_in3.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),       // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),      // reset_in3.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),       // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),      // reset_in3.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.reset_in1      (~ddr3_afi_reset_export_reset),       // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.reset_in3      (cpu_debug_reset_request_reset),      // reset_in3.reset
		.clk            (vga_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (ddr3_afi_clk_clk),                   //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
